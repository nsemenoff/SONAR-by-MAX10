
module main_clock (
	clkout,
	oscena);	

	output		clkout;
	input		oscena;
endmodule
